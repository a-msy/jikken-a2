/*
 * This code is produced by: 
 *   FSL Compiler version 0.1 alpha (2020-05-19) build 20E314
 *   Designed by Nobuya WATANABE, Okayama University, 2015-2020.
 * 
 *   Mon Jun 08 23:18:45 JST 2020
 * 
 * The source file of this code: 'mult32.fsl'.
 * 
 * INFO: 
 * 
 */
/* ModuleDef: mult32 */

module mult32(p_reset, m_clock, a, b, out, en, mult);
  input         p_reset;
  wire          p_reset;
  input         m_clock;
  wire          m_clock;
  input  [31:0] a;
  wire   [31:0] a;
  input  [31:0] b;
  wire   [31:0] b;
  output [63:0] out;
  wire   [63:0] out;
  output        en;
  wire          en;
  input         mult;
  wire          mult;
  /* for bundle-type input/output */
  /* local decls */
  wire          __net0;
  wire          __net1;
  wire          __net10;
  wire          __net11;
  wire          __net12;
  wire          __net13;
  wire          __net14;
  wire          __net15;
  wire          __net16;
  wire          __net17;
  wire          __net18;
  wire          __net19;
  wire          __net2;
  wire          __net20;
  wire          __net21;
  wire          __net22;
  wire          __net23;
  wire          __net24;
  wire          __net25;
  wire          __net26;
  wire          __net27;
  wire          __net28;
  wire          __net29;
  wire          __net3;
  wire          __net30;
  wire          __net31;
  wire   [63:0] __net32;
  wire          __net4;
  wire          __net5;
  wire          __net6;
  wire          __net7;
  wire          __net8;
  wire          __net9;
  /* assigns */
  assign __net0 = mult ? b[0:0] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net1 = mult ? b[1:1] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net10 = mult ? b[10:10] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net11 = mult ? b[11:11] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net12 = mult ? b[12:12] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net13 = mult ? b[13:13] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net14 = mult ? b[14:14] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net15 = mult ? b[15:15] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net16 = mult ? b[16:16] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net17 = mult ? b[17:17] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net18 = mult ? b[18:18] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net19 = mult ? b[19:19] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net2 = mult ? b[2:2] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net20 = mult ? b[20:20] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net21 = mult ? b[21:21] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net22 = mult ? b[22:22] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net23 = mult ? b[23:23] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net24 = mult ? b[24:24] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net25 = mult ? b[25:25] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net26 = mult ? b[26:26] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net27 = mult ? b[27:27] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net28 = mult ? b[28:28] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net29 = mult ? b[29:29] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net3 = mult ? b[3:3] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net30 = mult ? b[30:30] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net31 = mult ? b[31:31] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net32 = mult ? 
                     ((b[0:0] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 32) + ((b[1:1] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 31) + ((b[2:2] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 30) + ((b[3:3] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 29) + ((b[4:4] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 28) + ((b[5:5] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 27) + ((b[6:6] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 26) + ((b[7:7] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 25) + ((b[8:8] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 24) + ((b[9:9] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 23) + ((b[10:10] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 22) + ((b[11:11] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 21) + ((b[12:12] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 20) + ((b[13:13] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 19) + ((b[14:14] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 18) + ((b[15:15] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 17) + ((b[16:16] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 16) + ((b[17:17] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 15) + ((b[18:18] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 14) + ((b[19:19] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 13) + ((b[20:20] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 12) + ((b[21:21] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 11) + ((b[22:22] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 10) + ((b[23:23] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 9) + ((b[24:24] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 8) + ((b[25:25] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 7) + ((b[26:26] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 6) + ((b[27:27] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 5) + ((b[28:28] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 4) + ((b[29:29] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 3) + ((b[30:30] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 2) + ((b[31:31] == 1'B1 ? 
                       {a, 32'B00000000000000000000000000000000} : 
                       64'B0000000000000000000000000000000000000000000000000000000000000000) >> 1) : 
                     64'bx;
  assign __net4 = mult ? b[4:4] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net5 = mult ? b[5:5] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net6 = mult ? b[6:6] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net7 = mult ? b[7:7] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net8 = mult ? b[8:8] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign __net9 = mult ? b[9:9] == 1'B1 ? 1'b1 : 1'b0 : 1'bx;
  assign out = mult ? __net32 : 64'bx;
  /* invokes */
  /* private function */
  assign en = mult;
  /* defs */
  /* FunDef mult */
  /*   parameter: a: Bit(32) */
  /*   parameter: b: Bit(32) */
endmodule
/* End of file (mult32.v) */
